-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bb9",
     9 => x"90080b0b",
    10 => x"0bb99408",
    11 => x"0b0b0bb9",
    12 => x"98080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b9980c0b",
    16 => x"0b0bb994",
    17 => x"0c0b0b0b",
    18 => x"b9900c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb1fc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b9907080",
    57 => x"c3cc278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"51888804",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb9a00c",
    65 => x"9f0bb9a4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b9a408ff",
    69 => x"05b9a40c",
    70 => x"b9a40880",
    71 => x"25eb38b9",
    72 => x"a008ff05",
    73 => x"b9a00cb9",
    74 => x"a0088025",
    75 => x"d738800b",
    76 => x"b9a40c80",
    77 => x"0bb9a00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb9a008",
    97 => x"258f3882",
    98 => x"bd2db9a0",
    99 => x"08ff05b9",
   100 => x"a00c82ff",
   101 => x"04b9a008",
   102 => x"b9a40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b9a008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b9a4",
   111 => x"088105b9",
   112 => x"a40cb9a4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb9a40c",
   116 => x"b9a00881",
   117 => x"05b9a00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b9",
   122 => x"a4088105",
   123 => x"b9a40cb9",
   124 => x"a408a02e",
   125 => x"0981068e",
   126 => x"38800bb9",
   127 => x"a40cb9a0",
   128 => x"088105b9",
   129 => x"a00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb9a8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb9a80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b9",
   169 => x"a8088407",
   170 => x"b9a80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb5b4",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfecc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b9a80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b9900c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"8dab2d80",
   203 => x"518cde2d",
   204 => x"8cde2d8c",
   205 => x"de2d8cde",
   206 => x"2d70f00c",
   207 => x"70f40c70",
   208 => x"f80c8111",
   209 => x"51907125",
   210 => x"e4388d98",
   211 => x"2d028405",
   212 => x"0d0402fc",
   213 => x"050dec51",
   214 => x"83710c82",
   215 => x"710c0284",
   216 => x"050d0402",
   217 => x"dc050d80",
   218 => x"59810bec",
   219 => x"0c840bec",
   220 => x"0c7a52b9",
   221 => x"ac51a9a0",
   222 => x"2db99008",
   223 => x"792e80f9",
   224 => x"38b9b008",
   225 => x"79ff1256",
   226 => x"59567379",
   227 => x"2e8b3881",
   228 => x"1874812a",
   229 => x"555873f7",
   230 => x"38f71858",
   231 => x"81598076",
   232 => x"2580d038",
   233 => x"77527351",
   234 => x"848b2dba",
   235 => x"8452b9ac",
   236 => x"51abdf2d",
   237 => x"b9900880",
   238 => x"2e9a38ba",
   239 => x"845783fc",
   240 => x"55767084",
   241 => x"055808e8",
   242 => x"0cfc1555",
   243 => x"748025f1",
   244 => x"3887db04",
   245 => x"b9900859",
   246 => x"848056b9",
   247 => x"ac51abb1",
   248 => x"2dfc8016",
   249 => x"81155556",
   250 => x"758024ff",
   251 => x"b7387880",
   252 => x"2e8738b5",
   253 => x"b85187fc",
   254 => x"04b6e451",
   255 => x"8fa82d78",
   256 => x"b9900c02",
   257 => x"a4050d04",
   258 => x"02f4050d",
   259 => x"810bec0c",
   260 => x"8cf92d89",
   261 => x"c82d81f8",
   262 => x"2d83528c",
   263 => x"de2d8151",
   264 => x"84f02dff",
   265 => x"12527180",
   266 => x"25f13888",
   267 => x"0bb6b00b",
   268 => x"81b72d88",
   269 => x"0bb6bc0b",
   270 => x"81b72d88",
   271 => x"0bb6c80b",
   272 => x"81b72d84",
   273 => x"0bec0cb3",
   274 => x"c45185fe",
   275 => x"2da09f2d",
   276 => x"b9900880",
   277 => x"2e80dc38",
   278 => x"b3dc5185",
   279 => x"fe2db3f4",
   280 => x"5186e32d",
   281 => x"86e351b1",
   282 => x"f42d8d98",
   283 => x"2d89d42d",
   284 => x"8fb82db5",
   285 => x"cc0b80f5",
   286 => x"2db9e408",
   287 => x"81065353",
   288 => x"71802e85",
   289 => x"38728407",
   290 => x"5372fc0c",
   291 => x"b6b00b80",
   292 => x"f52df00c",
   293 => x"b6bc0b80",
   294 => x"f52df40c",
   295 => x"b6c80b80",
   296 => x"f52df80c",
   297 => x"8652b990",
   298 => x"08833884",
   299 => x"5271ec0c",
   300 => x"88ed0480",
   301 => x"0bb9900c",
   302 => x"028c050d",
   303 => x"0471980c",
   304 => x"04ffb008",
   305 => x"b9900c04",
   306 => x"810bffb0",
   307 => x"0c04800b",
   308 => x"ffb00c04",
   309 => x"02f4050d",
   310 => x"8ad604b9",
   311 => x"900881f0",
   312 => x"2e098106",
   313 => x"8938810b",
   314 => x"b7c80c8a",
   315 => x"d604b990",
   316 => x"0881e02e",
   317 => x"09810689",
   318 => x"38810bb7",
   319 => x"cc0c8ad6",
   320 => x"04b99008",
   321 => x"52b7cc08",
   322 => x"802e8838",
   323 => x"b9900881",
   324 => x"80055271",
   325 => x"842c728f",
   326 => x"065353b7",
   327 => x"c808802e",
   328 => x"99387284",
   329 => x"29b78805",
   330 => x"72138171",
   331 => x"2b700973",
   332 => x"0806730c",
   333 => x"5153538a",
   334 => x"cc047284",
   335 => x"29b78805",
   336 => x"72138371",
   337 => x"2b720807",
   338 => x"720c5353",
   339 => x"800bb7cc",
   340 => x"0c800bb7",
   341 => x"c80cb9b8",
   342 => x"518bd72d",
   343 => x"b99008ff",
   344 => x"24fef838",
   345 => x"800bb990",
   346 => x"0c028c05",
   347 => x"0d0402f8",
   348 => x"050db788",
   349 => x"528f5180",
   350 => x"72708405",
   351 => x"540cff11",
   352 => x"51708025",
   353 => x"f2380288",
   354 => x"050d0402",
   355 => x"f0050d75",
   356 => x"5189ce2d",
   357 => x"70822cfc",
   358 => x"06b78811",
   359 => x"72109e06",
   360 => x"71087072",
   361 => x"2a708306",
   362 => x"82742b70",
   363 => x"09740676",
   364 => x"0c545156",
   365 => x"57535153",
   366 => x"89c82d71",
   367 => x"b9900c02",
   368 => x"90050d04",
   369 => x"02fc050d",
   370 => x"72518071",
   371 => x"0c800b84",
   372 => x"120c0284",
   373 => x"050d0402",
   374 => x"f0050d75",
   375 => x"70088412",
   376 => x"08535353",
   377 => x"ff547171",
   378 => x"2ea83889",
   379 => x"ce2d8413",
   380 => x"08708429",
   381 => x"14881170",
   382 => x"087081ff",
   383 => x"06841808",
   384 => x"81118706",
   385 => x"841a0c53",
   386 => x"51555151",
   387 => x"5189c82d",
   388 => x"715473b9",
   389 => x"900c0290",
   390 => x"050d0402",
   391 => x"f8050d89",
   392 => x"ce2de008",
   393 => x"708b2a70",
   394 => x"81065152",
   395 => x"5270802e",
   396 => x"9d38b9b8",
   397 => x"08708429",
   398 => x"b9c00573",
   399 => x"81ff0671",
   400 => x"0c5151b9",
   401 => x"b8088111",
   402 => x"8706b9b8",
   403 => x"0c51800b",
   404 => x"b9e00c89",
   405 => x"c12d89c8",
   406 => x"2d028805",
   407 => x"0d0402fc",
   408 => x"050d89ce",
   409 => x"2d810bb9",
   410 => x"e00c89c8",
   411 => x"2db9e008",
   412 => x"5170fa38",
   413 => x"0284050d",
   414 => x"0402fc05",
   415 => x"0db9b851",
   416 => x"8bc42d8a",
   417 => x"ee2d8c9b",
   418 => x"5189bd2d",
   419 => x"0284050d",
   420 => x"04b9f008",
   421 => x"b9900c04",
   422 => x"02fc050d",
   423 => x"810bb7d0",
   424 => x"0c815184",
   425 => x"f02d0284",
   426 => x"050d0402",
   427 => x"fc050d8d",
   428 => x"b50489d4",
   429 => x"2d80f851",
   430 => x"8b8b2db9",
   431 => x"9008f338",
   432 => x"80da518b",
   433 => x"8b2db990",
   434 => x"08e838b9",
   435 => x"9008b7d0",
   436 => x"0cb99008",
   437 => x"5184f02d",
   438 => x"0284050d",
   439 => x"0402ec05",
   440 => x"0d765480",
   441 => x"52870b88",
   442 => x"1580f52d",
   443 => x"56537472",
   444 => x"248338a0",
   445 => x"53725182",
   446 => x"f92d8112",
   447 => x"8b1580f5",
   448 => x"2d545272",
   449 => x"7225de38",
   450 => x"0294050d",
   451 => x"0402f005",
   452 => x"0db9f008",
   453 => x"5481f82d",
   454 => x"800bb9f4",
   455 => x"0c730880",
   456 => x"2e818038",
   457 => x"820bb9a4",
   458 => x"0cb9f408",
   459 => x"8f06b9a0",
   460 => x"0c730852",
   461 => x"71832e96",
   462 => x"38718326",
   463 => x"89387181",
   464 => x"2eaf388f",
   465 => x"8e047185",
   466 => x"2e9f388f",
   467 => x"8e048814",
   468 => x"80f52d84",
   469 => x"1508b480",
   470 => x"53545285",
   471 => x"fe2d7184",
   472 => x"29137008",
   473 => x"52528f92",
   474 => x"0473518d",
   475 => x"dd2d8f8e",
   476 => x"04b9e408",
   477 => x"8815082c",
   478 => x"70810651",
   479 => x"5271802e",
   480 => x"8738b484",
   481 => x"518f8b04",
   482 => x"b4885185",
   483 => x"fe2d8414",
   484 => x"085185fe",
   485 => x"2db9f408",
   486 => x"8105b9f4",
   487 => x"0c8c1454",
   488 => x"8e9d0402",
   489 => x"90050d04",
   490 => x"71b9f00c",
   491 => x"8e8d2db9",
   492 => x"f408ff05",
   493 => x"b9f80c04",
   494 => x"02e8050d",
   495 => x"b9f008b9",
   496 => x"fc085755",
   497 => x"80f8518b",
   498 => x"8b2db990",
   499 => x"08812a70",
   500 => x"81065152",
   501 => x"71802ea1",
   502 => x"388fdf04",
   503 => x"89d42d80",
   504 => x"f8518b8b",
   505 => x"2db99008",
   506 => x"f338b7d0",
   507 => x"08813270",
   508 => x"b7d00c70",
   509 => x"525284f0",
   510 => x"2d800bb9",
   511 => x"e80c800b",
   512 => x"b9ec0cb7",
   513 => x"d00882dd",
   514 => x"3880da51",
   515 => x"8b8b2db9",
   516 => x"9008802e",
   517 => x"8a38b9e8",
   518 => x"08818007",
   519 => x"b9e80c80",
   520 => x"d9518b8b",
   521 => x"2db99008",
   522 => x"802e8a38",
   523 => x"b9e80880",
   524 => x"c007b9e8",
   525 => x"0c819451",
   526 => x"8b8b2db9",
   527 => x"9008802e",
   528 => x"8938b9e8",
   529 => x"089007b9",
   530 => x"e80c8191",
   531 => x"518b8b2d",
   532 => x"b9900880",
   533 => x"2e8938b9",
   534 => x"e808a007",
   535 => x"b9e80c81",
   536 => x"f5518b8b",
   537 => x"2db99008",
   538 => x"802e8938",
   539 => x"b9e80881",
   540 => x"07b9e80c",
   541 => x"81f2518b",
   542 => x"8b2db990",
   543 => x"08802e89",
   544 => x"38b9e808",
   545 => x"8207b9e8",
   546 => x"0c81eb51",
   547 => x"8b8b2db9",
   548 => x"9008802e",
   549 => x"8938b9e8",
   550 => x"088407b9",
   551 => x"e80c81f4",
   552 => x"518b8b2d",
   553 => x"b9900880",
   554 => x"2e8938b9",
   555 => x"e8088807",
   556 => x"b9e80c80",
   557 => x"d8518b8b",
   558 => x"2db99008",
   559 => x"802e8a38",
   560 => x"b9ec0881",
   561 => x"8007b9ec",
   562 => x"0c92518b",
   563 => x"8b2db990",
   564 => x"08802e8a",
   565 => x"38b9ec08",
   566 => x"80c007b9",
   567 => x"ec0c9451",
   568 => x"8b8b2db9",
   569 => x"9008802e",
   570 => x"8938b9ec",
   571 => x"089007b9",
   572 => x"ec0c9151",
   573 => x"8b8b2db9",
   574 => x"9008802e",
   575 => x"8938b9ec",
   576 => x"08a007b9",
   577 => x"ec0c9d51",
   578 => x"8b8b2db9",
   579 => x"9008802e",
   580 => x"8938b9ec",
   581 => x"088107b9",
   582 => x"ec0c9b51",
   583 => x"8b8b2db9",
   584 => x"9008802e",
   585 => x"8938b9ec",
   586 => x"088207b9",
   587 => x"ec0c9c51",
   588 => x"8b8b2db9",
   589 => x"9008802e",
   590 => x"8938b9ec",
   591 => x"088407b9",
   592 => x"ec0ca351",
   593 => x"8b8b2db9",
   594 => x"9008802e",
   595 => x"8938b9ec",
   596 => x"088807b9",
   597 => x"ec0c81fd",
   598 => x"518b8b2d",
   599 => x"81fa518b",
   600 => x"8b2d9896",
   601 => x"0481f551",
   602 => x"8b8b2db9",
   603 => x"9008812a",
   604 => x"70810651",
   605 => x"5271802e",
   606 => x"af38b9f8",
   607 => x"08527180",
   608 => x"2e8938ff",
   609 => x"12b9f80c",
   610 => x"93a804b9",
   611 => x"f40810b9",
   612 => x"f4080570",
   613 => x"84291651",
   614 => x"52881208",
   615 => x"802e8938",
   616 => x"ff518812",
   617 => x"0852712d",
   618 => x"81f2518b",
   619 => x"8b2db990",
   620 => x"08812a70",
   621 => x"81065152",
   622 => x"71802eb1",
   623 => x"38b9f408",
   624 => x"ff11b9f8",
   625 => x"08565353",
   626 => x"73722589",
   627 => x"388114b9",
   628 => x"f80c93ed",
   629 => x"04721013",
   630 => x"70842916",
   631 => x"51528812",
   632 => x"08802e89",
   633 => x"38fe5188",
   634 => x"12085271",
   635 => x"2d81fd51",
   636 => x"8b8b2db9",
   637 => x"9008812a",
   638 => x"70810651",
   639 => x"5271802e",
   640 => x"ad38b9f8",
   641 => x"08802e89",
   642 => x"38800bb9",
   643 => x"f80c94ae",
   644 => x"04b9f408",
   645 => x"10b9f408",
   646 => x"05708429",
   647 => x"16515288",
   648 => x"1208802e",
   649 => x"8938fd51",
   650 => x"88120852",
   651 => x"712d81fa",
   652 => x"518b8b2d",
   653 => x"b9900881",
   654 => x"2a708106",
   655 => x"51527180",
   656 => x"2eae38b9",
   657 => x"f408ff11",
   658 => x"5452b9f8",
   659 => x"08732588",
   660 => x"3872b9f8",
   661 => x"0c94f004",
   662 => x"71101270",
   663 => x"84291651",
   664 => x"52881208",
   665 => x"802e8938",
   666 => x"fc518812",
   667 => x"0852712d",
   668 => x"b9f80870",
   669 => x"53547380",
   670 => x"2e8a388c",
   671 => x"15ff1555",
   672 => x"5594f604",
   673 => x"820bb9a4",
   674 => x"0c718f06",
   675 => x"b9a00c81",
   676 => x"eb518b8b",
   677 => x"2db99008",
   678 => x"812a7081",
   679 => x"06515271",
   680 => x"802ead38",
   681 => x"7408852e",
   682 => x"098106a4",
   683 => x"38881580",
   684 => x"f52dff05",
   685 => x"52718816",
   686 => x"81b72d71",
   687 => x"982b5271",
   688 => x"80258838",
   689 => x"800b8816",
   690 => x"81b72d74",
   691 => x"518ddd2d",
   692 => x"81f4518b",
   693 => x"8b2db990",
   694 => x"08812a70",
   695 => x"81065152",
   696 => x"71802eb3",
   697 => x"38740885",
   698 => x"2e098106",
   699 => x"aa388815",
   700 => x"80f52d81",
   701 => x"05527188",
   702 => x"1681b72d",
   703 => x"7181ff06",
   704 => x"8b1680f5",
   705 => x"2d545272",
   706 => x"72278738",
   707 => x"72881681",
   708 => x"b72d7451",
   709 => x"8ddd2d80",
   710 => x"da518b8b",
   711 => x"2db99008",
   712 => x"812a7081",
   713 => x"06515271",
   714 => x"802e81a6",
   715 => x"38b9f008",
   716 => x"b9f80855",
   717 => x"5373802e",
   718 => x"8a388c13",
   719 => x"ff155553",
   720 => x"96b50472",
   721 => x"08527182",
   722 => x"2ea63871",
   723 => x"82268938",
   724 => x"71812ea9",
   725 => x"3897d204",
   726 => x"71832eb1",
   727 => x"3871842e",
   728 => x"09810680",
   729 => x"ed388813",
   730 => x"08518fa8",
   731 => x"2d97d204",
   732 => x"b9f80851",
   733 => x"88130852",
   734 => x"712d97d2",
   735 => x"04810b88",
   736 => x"14082bb9",
   737 => x"e40832b9",
   738 => x"e40c97a8",
   739 => x"04881380",
   740 => x"f52d8105",
   741 => x"8b1480f5",
   742 => x"2d535471",
   743 => x"74248338",
   744 => x"80547388",
   745 => x"1481b72d",
   746 => x"8e8d2d97",
   747 => x"d2047508",
   748 => x"802ea238",
   749 => x"7508518b",
   750 => x"8b2db990",
   751 => x"08810652",
   752 => x"71802e8b",
   753 => x"38b9f808",
   754 => x"51841608",
   755 => x"52712d88",
   756 => x"165675da",
   757 => x"38805480",
   758 => x"0bb9a40c",
   759 => x"738f06b9",
   760 => x"a00ca052",
   761 => x"73b9f808",
   762 => x"2e098106",
   763 => x"9838b9f4",
   764 => x"08ff0574",
   765 => x"32700981",
   766 => x"05707207",
   767 => x"9f2a9171",
   768 => x"31515153",
   769 => x"53715182",
   770 => x"f92d8114",
   771 => x"548e7425",
   772 => x"c638b7d0",
   773 => x"085271b9",
   774 => x"900c0298",
   775 => x"050d0402",
   776 => x"f4050dd4",
   777 => x"5281ff72",
   778 => x"0c710853",
   779 => x"81ff720c",
   780 => x"72882b83",
   781 => x"fe800672",
   782 => x"087081ff",
   783 => x"06515253",
   784 => x"81ff720c",
   785 => x"72710788",
   786 => x"2b720870",
   787 => x"81ff0651",
   788 => x"525381ff",
   789 => x"720c7271",
   790 => x"07882b72",
   791 => x"087081ff",
   792 => x"067207b9",
   793 => x"900c5253",
   794 => x"028c050d",
   795 => x"0402f405",
   796 => x"0d747671",
   797 => x"81ff06d4",
   798 => x"0c5353ba",
   799 => x"80088538",
   800 => x"71892b52",
   801 => x"71982ad4",
   802 => x"0c71902a",
   803 => x"7081ff06",
   804 => x"d40c5171",
   805 => x"882a7081",
   806 => x"ff06d40c",
   807 => x"517181ff",
   808 => x"06d40c72",
   809 => x"902a7081",
   810 => x"ff06d40c",
   811 => x"51d40870",
   812 => x"81ff0651",
   813 => x"5182b8bf",
   814 => x"527081ff",
   815 => x"2e098106",
   816 => x"943881ff",
   817 => x"0bd40cd4",
   818 => x"087081ff",
   819 => x"06ff1454",
   820 => x"515171e5",
   821 => x"3870b990",
   822 => x"0c028c05",
   823 => x"0d0402fc",
   824 => x"050d81c7",
   825 => x"5181ff0b",
   826 => x"d40cff11",
   827 => x"51708025",
   828 => x"f4380284",
   829 => x"050d0402",
   830 => x"f4050d81",
   831 => x"ff0bd40c",
   832 => x"93538052",
   833 => x"87fc80c1",
   834 => x"5198ed2d",
   835 => x"b990088b",
   836 => x"3881ff0b",
   837 => x"d40c8153",
   838 => x"9aa40499",
   839 => x"de2dff13",
   840 => x"5372df38",
   841 => x"72b9900c",
   842 => x"028c050d",
   843 => x"0402ec05",
   844 => x"0d810bba",
   845 => x"800c8454",
   846 => x"d008708f",
   847 => x"2a708106",
   848 => x"51515372",
   849 => x"f33872d0",
   850 => x"0c99de2d",
   851 => x"b48c5185",
   852 => x"fe2dd008",
   853 => x"708f2a70",
   854 => x"81065151",
   855 => x"5372f338",
   856 => x"810bd00c",
   857 => x"b1538052",
   858 => x"84d480c0",
   859 => x"5198ed2d",
   860 => x"b9900881",
   861 => x"2e933872",
   862 => x"822ebd38",
   863 => x"ff135372",
   864 => x"e538ff14",
   865 => x"5473ffb0",
   866 => x"3899de2d",
   867 => x"83aa5284",
   868 => x"9c80c851",
   869 => x"98ed2db9",
   870 => x"9008812e",
   871 => x"09810692",
   872 => x"38989f2d",
   873 => x"b9900883",
   874 => x"ffff0653",
   875 => x"7283aa2e",
   876 => x"9d3899f7",
   877 => x"2d9bc904",
   878 => x"b4985185",
   879 => x"fe2d8053",
   880 => x"9d9704b4",
   881 => x"b05185fe",
   882 => x"2d80549c",
   883 => x"e90481ff",
   884 => x"0bd40cb1",
   885 => x"5499de2d",
   886 => x"8fcf5380",
   887 => x"5287fc80",
   888 => x"f75198ed",
   889 => x"2db99008",
   890 => x"55b99008",
   891 => x"812e0981",
   892 => x"069b3881",
   893 => x"ff0bd40c",
   894 => x"820a5284",
   895 => x"9c80e951",
   896 => x"98ed2db9",
   897 => x"9008802e",
   898 => x"8d3899de",
   899 => x"2dff1353",
   900 => x"72c9389c",
   901 => x"dc0481ff",
   902 => x"0bd40cb9",
   903 => x"90085287",
   904 => x"fc80fa51",
   905 => x"98ed2db9",
   906 => x"9008b138",
   907 => x"81ff0bd4",
   908 => x"0cd40853",
   909 => x"81ff0bd4",
   910 => x"0c81ff0b",
   911 => x"d40c81ff",
   912 => x"0bd40c81",
   913 => x"ff0bd40c",
   914 => x"72862a70",
   915 => x"81067656",
   916 => x"51537295",
   917 => x"38b99008",
   918 => x"549ce904",
   919 => x"73822efe",
   920 => x"e238ff14",
   921 => x"5473feed",
   922 => x"3873ba80",
   923 => x"0c738b38",
   924 => x"815287fc",
   925 => x"80d05198",
   926 => x"ed2d81ff",
   927 => x"0bd40cd0",
   928 => x"08708f2a",
   929 => x"70810651",
   930 => x"515372f3",
   931 => x"3872d00c",
   932 => x"81ff0bd4",
   933 => x"0c815372",
   934 => x"b9900c02",
   935 => x"94050d04",
   936 => x"02e8050d",
   937 => x"78558056",
   938 => x"81ff0bd4",
   939 => x"0cd00870",
   940 => x"8f2a7081",
   941 => x"06515153",
   942 => x"72f33882",
   943 => x"810bd00c",
   944 => x"81ff0bd4",
   945 => x"0c775287",
   946 => x"fc80d151",
   947 => x"98ed2d80",
   948 => x"dbc6df54",
   949 => x"b9900880",
   950 => x"2e8a38b4",
   951 => x"d05185fe",
   952 => x"2d9eb704",
   953 => x"81ff0bd4",
   954 => x"0cd40870",
   955 => x"81ff0651",
   956 => x"537281fe",
   957 => x"2e098106",
   958 => x"9d3880ff",
   959 => x"53989f2d",
   960 => x"b9900875",
   961 => x"70840557",
   962 => x"0cff1353",
   963 => x"728025ed",
   964 => x"3881569e",
   965 => x"9c04ff14",
   966 => x"5473c938",
   967 => x"81ff0bd4",
   968 => x"0c81ff0b",
   969 => x"d40cd008",
   970 => x"708f2a70",
   971 => x"81065151",
   972 => x"5372f338",
   973 => x"72d00c75",
   974 => x"b9900c02",
   975 => x"98050d04",
   976 => x"02e8050d",
   977 => x"77797b58",
   978 => x"55558053",
   979 => x"727625a3",
   980 => x"38747081",
   981 => x"055680f5",
   982 => x"2d747081",
   983 => x"055680f5",
   984 => x"2d525271",
   985 => x"712e8638",
   986 => x"81519ef5",
   987 => x"04811353",
   988 => x"9ecc0480",
   989 => x"5170b990",
   990 => x"0c029805",
   991 => x"0d0402ec",
   992 => x"050d7655",
   993 => x"74802ebe",
   994 => x"389a1580",
   995 => x"e02d51ac",
   996 => x"b82db990",
   997 => x"08b99008",
   998 => x"80c0b40c",
   999 => x"b9900854",
  1000 => x"5480c090",
  1001 => x"08802e99",
  1002 => x"38941580",
  1003 => x"e02d51ac",
  1004 => x"b82db990",
  1005 => x"08902b83",
  1006 => x"fff00a06",
  1007 => x"70750751",
  1008 => x"537280c0",
  1009 => x"b40c80c0",
  1010 => x"b4085372",
  1011 => x"802e9d38",
  1012 => x"80c08808",
  1013 => x"fe147129",
  1014 => x"80c09c08",
  1015 => x"0580c0b8",
  1016 => x"0c70842b",
  1017 => x"80c0940c",
  1018 => x"54a09a04",
  1019 => x"80c0a008",
  1020 => x"80c0b40c",
  1021 => x"80c0a408",
  1022 => x"80c0b80c",
  1023 => x"80c09008",
  1024 => x"802e8b38",
  1025 => x"80c08808",
  1026 => x"842b53a0",
  1027 => x"950480c0",
  1028 => x"a808842b",
  1029 => x"537280c0",
  1030 => x"940c0294",
  1031 => x"050d0402",
  1032 => x"d8050d80",
  1033 => x"0b80c090",
  1034 => x"0c84549a",
  1035 => x"ad2db990",
  1036 => x"08802e95",
  1037 => x"38ba8452",
  1038 => x"80519da0",
  1039 => x"2db99008",
  1040 => x"802e8638",
  1041 => x"fe54a0d1",
  1042 => x"04ff1454",
  1043 => x"738024db",
  1044 => x"38738c38",
  1045 => x"b4e05185",
  1046 => x"fe2d7355",
  1047 => x"a5f30480",
  1048 => x"56810b80",
  1049 => x"c0bc0c88",
  1050 => x"53b4f452",
  1051 => x"baba519e",
  1052 => x"c02db990",
  1053 => x"08762e09",
  1054 => x"81068838",
  1055 => x"b9900880",
  1056 => x"c0bc0c88",
  1057 => x"53b58052",
  1058 => x"bad6519e",
  1059 => x"c02db990",
  1060 => x"088838b9",
  1061 => x"900880c0",
  1062 => x"bc0c80c0",
  1063 => x"bc08802e",
  1064 => x"80f638bd",
  1065 => x"ca0b80f5",
  1066 => x"2dbdcb0b",
  1067 => x"80f52d71",
  1068 => x"982b7190",
  1069 => x"2b07bdcc",
  1070 => x"0b80f52d",
  1071 => x"70882b72",
  1072 => x"07bdcd0b",
  1073 => x"80f52d71",
  1074 => x"07be820b",
  1075 => x"80f52dbe",
  1076 => x"830b80f5",
  1077 => x"2d71882b",
  1078 => x"07535f54",
  1079 => x"525a5657",
  1080 => x"557381ab",
  1081 => x"aa2e0981",
  1082 => x"068d3875",
  1083 => x"51ac882d",
  1084 => x"b9900856",
  1085 => x"a2840473",
  1086 => x"82d4d52e",
  1087 => x"8738b58c",
  1088 => x"51a2c604",
  1089 => x"ba845275",
  1090 => x"519da02d",
  1091 => x"b9900855",
  1092 => x"b9900880",
  1093 => x"2e83dc38",
  1094 => x"8853b580",
  1095 => x"52bad651",
  1096 => x"9ec02db9",
  1097 => x"90088a38",
  1098 => x"810b80c0",
  1099 => x"900ca2cc",
  1100 => x"048853b4",
  1101 => x"f452baba",
  1102 => x"519ec02d",
  1103 => x"b9900880",
  1104 => x"2e8a38b5",
  1105 => x"a05185fe",
  1106 => x"2da3a604",
  1107 => x"be820b80",
  1108 => x"f52d5473",
  1109 => x"80d52e09",
  1110 => x"810680ca",
  1111 => x"38be830b",
  1112 => x"80f52d54",
  1113 => x"7381aa2e",
  1114 => x"098106ba",
  1115 => x"38800bba",
  1116 => x"840b80f5",
  1117 => x"2d565474",
  1118 => x"81e92e83",
  1119 => x"38815474",
  1120 => x"81eb2e8c",
  1121 => x"38805573",
  1122 => x"752e0981",
  1123 => x"0682e438",
  1124 => x"ba8f0b80",
  1125 => x"f52d5574",
  1126 => x"8d38ba90",
  1127 => x"0b80f52d",
  1128 => x"5473822e",
  1129 => x"86388055",
  1130 => x"a5f304ba",
  1131 => x"910b80f5",
  1132 => x"2d7080c0",
  1133 => x"880cff05",
  1134 => x"80c08c0c",
  1135 => x"ba920b80",
  1136 => x"f52dba93",
  1137 => x"0b80f52d",
  1138 => x"58760577",
  1139 => x"82802905",
  1140 => x"7080c098",
  1141 => x"0cba940b",
  1142 => x"80f52d70",
  1143 => x"80c0ac0c",
  1144 => x"80c09008",
  1145 => x"59575876",
  1146 => x"802e81ac",
  1147 => x"388853b5",
  1148 => x"8052bad6",
  1149 => x"519ec02d",
  1150 => x"b9900881",
  1151 => x"f63880c0",
  1152 => x"88087084",
  1153 => x"2b80c094",
  1154 => x"0c7080c0",
  1155 => x"a80cbaa9",
  1156 => x"0b80f52d",
  1157 => x"baa80b80",
  1158 => x"f52d7182",
  1159 => x"802905ba",
  1160 => x"aa0b80f5",
  1161 => x"2d708480",
  1162 => x"802912ba",
  1163 => x"ab0b80f5",
  1164 => x"2d708180",
  1165 => x"0a291270",
  1166 => x"80c0b00c",
  1167 => x"80c0ac08",
  1168 => x"712980c0",
  1169 => x"98080570",
  1170 => x"80c09c0c",
  1171 => x"bab10b80",
  1172 => x"f52dbab0",
  1173 => x"0b80f52d",
  1174 => x"71828029",
  1175 => x"05bab20b",
  1176 => x"80f52d70",
  1177 => x"84808029",
  1178 => x"12bab30b",
  1179 => x"80f52d70",
  1180 => x"982b81f0",
  1181 => x"0a067205",
  1182 => x"7080c0a0",
  1183 => x"0cfe117e",
  1184 => x"29770580",
  1185 => x"c0a40c52",
  1186 => x"59524354",
  1187 => x"5e515259",
  1188 => x"525d5759",
  1189 => x"57a5ec04",
  1190 => x"ba960b80",
  1191 => x"f52dba95",
  1192 => x"0b80f52d",
  1193 => x"71828029",
  1194 => x"057080c0",
  1195 => x"940c70a0",
  1196 => x"2983ff05",
  1197 => x"70892a70",
  1198 => x"80c0a80c",
  1199 => x"ba9b0b80",
  1200 => x"f52dba9a",
  1201 => x"0b80f52d",
  1202 => x"71828029",
  1203 => x"057080c0",
  1204 => x"b00c7b71",
  1205 => x"291e7080",
  1206 => x"c0a40c7d",
  1207 => x"80c0a00c",
  1208 => x"730580c0",
  1209 => x"9c0c555e",
  1210 => x"51515555",
  1211 => x"80519efe",
  1212 => x"2d815574",
  1213 => x"b9900c02",
  1214 => x"a8050d04",
  1215 => x"02ec050d",
  1216 => x"7670872c",
  1217 => x"7180ff06",
  1218 => x"55565480",
  1219 => x"c090088a",
  1220 => x"3873882c",
  1221 => x"7481ff06",
  1222 => x"5455ba84",
  1223 => x"5280c098",
  1224 => x"0815519d",
  1225 => x"a02db990",
  1226 => x"0854b990",
  1227 => x"08802eb4",
  1228 => x"3880c090",
  1229 => x"08802e98",
  1230 => x"38728429",
  1231 => x"ba840570",
  1232 => x"085253ac",
  1233 => x"882db990",
  1234 => x"08f00a06",
  1235 => x"53a6e204",
  1236 => x"7210ba84",
  1237 => x"057080e0",
  1238 => x"2d5253ac",
  1239 => x"b82db990",
  1240 => x"08537254",
  1241 => x"73b9900c",
  1242 => x"0294050d",
  1243 => x"0402e005",
  1244 => x"0d797084",
  1245 => x"2c80c0b8",
  1246 => x"0805718f",
  1247 => x"06525553",
  1248 => x"728938ba",
  1249 => x"84527351",
  1250 => x"9da02d72",
  1251 => x"a029ba84",
  1252 => x"05548074",
  1253 => x"80f52d56",
  1254 => x"5374732e",
  1255 => x"83388153",
  1256 => x"7481e52e",
  1257 => x"81ef3881",
  1258 => x"70740654",
  1259 => x"5872802e",
  1260 => x"81e3388b",
  1261 => x"1480f52d",
  1262 => x"70832a79",
  1263 => x"06585676",
  1264 => x"9838b7d4",
  1265 => x"08537288",
  1266 => x"3872be84",
  1267 => x"0b81b72d",
  1268 => x"76b7d40c",
  1269 => x"7353a997",
  1270 => x"04758f2e",
  1271 => x"09810681",
  1272 => x"b438749f",
  1273 => x"068d29bd",
  1274 => x"f7115153",
  1275 => x"811480f5",
  1276 => x"2d737081",
  1277 => x"055581b7",
  1278 => x"2d831480",
  1279 => x"f52d7370",
  1280 => x"81055581",
  1281 => x"b72d8514",
  1282 => x"80f52d73",
  1283 => x"70810555",
  1284 => x"81b72d87",
  1285 => x"1480f52d",
  1286 => x"73708105",
  1287 => x"5581b72d",
  1288 => x"891480f5",
  1289 => x"2d737081",
  1290 => x"055581b7",
  1291 => x"2d8e1480",
  1292 => x"f52d7370",
  1293 => x"81055581",
  1294 => x"b72d9014",
  1295 => x"80f52d73",
  1296 => x"70810555",
  1297 => x"81b72d92",
  1298 => x"1480f52d",
  1299 => x"73708105",
  1300 => x"5581b72d",
  1301 => x"941480f5",
  1302 => x"2d737081",
  1303 => x"055581b7",
  1304 => x"2d961480",
  1305 => x"f52d7370",
  1306 => x"81055581",
  1307 => x"b72d9814",
  1308 => x"80f52d73",
  1309 => x"70810555",
  1310 => x"81b72d9c",
  1311 => x"1480f52d",
  1312 => x"73708105",
  1313 => x"5581b72d",
  1314 => x"9e1480f5",
  1315 => x"2d7381b7",
  1316 => x"2d77b7d4",
  1317 => x"0c805372",
  1318 => x"b9900c02",
  1319 => x"a0050d04",
  1320 => x"02cc050d",
  1321 => x"7e605e5a",
  1322 => x"800b80c0",
  1323 => x"b40880c0",
  1324 => x"b808595c",
  1325 => x"56805880",
  1326 => x"c0940878",
  1327 => x"2e81b038",
  1328 => x"778f06a0",
  1329 => x"17575473",
  1330 => x"8f38ba84",
  1331 => x"52765181",
  1332 => x"17579da0",
  1333 => x"2dba8456",
  1334 => x"807680f5",
  1335 => x"2d565474",
  1336 => x"742e8338",
  1337 => x"81547481",
  1338 => x"e52e80f7",
  1339 => x"38817075",
  1340 => x"06555c73",
  1341 => x"802e80eb",
  1342 => x"388b1680",
  1343 => x"f52d9806",
  1344 => x"597880df",
  1345 => x"388b537c",
  1346 => x"5275519e",
  1347 => x"c02db990",
  1348 => x"0880d038",
  1349 => x"9c160851",
  1350 => x"ac882db9",
  1351 => x"9008841b",
  1352 => x"0c9a1680",
  1353 => x"e02d51ac",
  1354 => x"b82db990",
  1355 => x"08b99008",
  1356 => x"881c0cb9",
  1357 => x"90085555",
  1358 => x"80c09008",
  1359 => x"802e9838",
  1360 => x"941680e0",
  1361 => x"2d51acb8",
  1362 => x"2db99008",
  1363 => x"902b83ff",
  1364 => x"f00a0670",
  1365 => x"16515473",
  1366 => x"881b0c78",
  1367 => x"7a0c7b54",
  1368 => x"aba80481",
  1369 => x"185880c0",
  1370 => x"94087826",
  1371 => x"fed23880",
  1372 => x"c0900880",
  1373 => x"2eb0387a",
  1374 => x"51a5fc2d",
  1375 => x"b99008b9",
  1376 => x"900880ff",
  1377 => x"fffff806",
  1378 => x"555b7380",
  1379 => x"fffffff8",
  1380 => x"2e9438b9",
  1381 => x"9008fe05",
  1382 => x"80c08808",
  1383 => x"2980c09c",
  1384 => x"080557a9",
  1385 => x"b5048054",
  1386 => x"73b9900c",
  1387 => x"02b4050d",
  1388 => x"0402f405",
  1389 => x"0d747008",
  1390 => x"8105710c",
  1391 => x"700880c0",
  1392 => x"8c080653",
  1393 => x"53718e38",
  1394 => x"88130851",
  1395 => x"a5fc2db9",
  1396 => x"90088814",
  1397 => x"0c810bb9",
  1398 => x"900c028c",
  1399 => x"050d0402",
  1400 => x"f0050d75",
  1401 => x"881108fe",
  1402 => x"0580c088",
  1403 => x"082980c0",
  1404 => x"9c081172",
  1405 => x"0880c08c",
  1406 => x"08060579",
  1407 => x"55535454",
  1408 => x"9da02d02",
  1409 => x"90050d04",
  1410 => x"02f4050d",
  1411 => x"7470882a",
  1412 => x"83fe8006",
  1413 => x"7072982a",
  1414 => x"0772882b",
  1415 => x"87fc8080",
  1416 => x"0673982b",
  1417 => x"81f00a06",
  1418 => x"71730707",
  1419 => x"b9900c56",
  1420 => x"51535102",
  1421 => x"8c050d04",
  1422 => x"02f8050d",
  1423 => x"028e0580",
  1424 => x"f52d7488",
  1425 => x"2b077083",
  1426 => x"ffff06b9",
  1427 => x"900c5102",
  1428 => x"88050d04",
  1429 => x"02f4050d",
  1430 => x"74767853",
  1431 => x"54528071",
  1432 => x"25973872",
  1433 => x"70810554",
  1434 => x"80f52d72",
  1435 => x"70810554",
  1436 => x"81b72dff",
  1437 => x"115170eb",
  1438 => x"38807281",
  1439 => x"b72d028c",
  1440 => x"050d0402",
  1441 => x"e8050d77",
  1442 => x"56807056",
  1443 => x"54737624",
  1444 => x"b33880c0",
  1445 => x"9408742e",
  1446 => x"ab387351",
  1447 => x"a6ed2db9",
  1448 => x"9008b990",
  1449 => x"08098105",
  1450 => x"70b99008",
  1451 => x"079f2a77",
  1452 => x"05811757",
  1453 => x"57535374",
  1454 => x"76248938",
  1455 => x"80c09408",
  1456 => x"7426d738",
  1457 => x"72b9900c",
  1458 => x"0298050d",
  1459 => x"0402f005",
  1460 => x"0db98c08",
  1461 => x"1651ad83",
  1462 => x"2db99008",
  1463 => x"802e9c38",
  1464 => x"8b53b990",
  1465 => x"0852be84",
  1466 => x"51acd42d",
  1467 => x"80c0c008",
  1468 => x"5473802e",
  1469 => x"8638be84",
  1470 => x"51732d02",
  1471 => x"90050d04",
  1472 => x"02dc050d",
  1473 => x"80705a55",
  1474 => x"74b98c08",
  1475 => x"25b13880",
  1476 => x"c0940875",
  1477 => x"2ea93878",
  1478 => x"51a6ed2d",
  1479 => x"b9900809",
  1480 => x"810570b9",
  1481 => x"9008079f",
  1482 => x"2a760581",
  1483 => x"1b5b5654",
  1484 => x"74b98c08",
  1485 => x"25893880",
  1486 => x"c0940879",
  1487 => x"26d93880",
  1488 => x"557880c0",
  1489 => x"94082781",
  1490 => x"d1387851",
  1491 => x"a6ed2db9",
  1492 => x"9008802e",
  1493 => x"81a538b9",
  1494 => x"90088b05",
  1495 => x"80f52d70",
  1496 => x"842a7081",
  1497 => x"06771078",
  1498 => x"842bbe84",
  1499 => x"0b80f52d",
  1500 => x"5c5c5351",
  1501 => x"55567380",
  1502 => x"2e80c838",
  1503 => x"7416822b",
  1504 => x"b0be0bb7",
  1505 => x"e0120c54",
  1506 => x"77753110",
  1507 => x"80c0c411",
  1508 => x"55569074",
  1509 => x"70810556",
  1510 => x"81b72da0",
  1511 => x"7481b72d",
  1512 => x"7681ff06",
  1513 => x"81165854",
  1514 => x"73802e89",
  1515 => x"389c53be",
  1516 => x"8452afbb",
  1517 => x"048b53b9",
  1518 => x"90085280",
  1519 => x"c0c61651",
  1520 => x"aff30474",
  1521 => x"16822bad",
  1522 => x"cd0bb7e0",
  1523 => x"120c5476",
  1524 => x"81ff0681",
  1525 => x"16585473",
  1526 => x"802e8938",
  1527 => x"9c53be84",
  1528 => x"52afea04",
  1529 => x"8b53b990",
  1530 => x"08527775",
  1531 => x"311080c0",
  1532 => x"c4055176",
  1533 => x"55acd42d",
  1534 => x"b08f0474",
  1535 => x"90297531",
  1536 => x"701080c0",
  1537 => x"c4055154",
  1538 => x"b9900874",
  1539 => x"81b72d81",
  1540 => x"1959748b",
  1541 => x"24a338ae",
  1542 => x"c1047490",
  1543 => x"29753170",
  1544 => x"1080c0c4",
  1545 => x"058c7731",
  1546 => x"57515480",
  1547 => x"7481b72d",
  1548 => x"9e14ff16",
  1549 => x"565474f3",
  1550 => x"3802a405",
  1551 => x"0d0402fc",
  1552 => x"050db98c",
  1553 => x"081351ad",
  1554 => x"832db990",
  1555 => x"08802e88",
  1556 => x"38b99008",
  1557 => x"519efe2d",
  1558 => x"800bb98c",
  1559 => x"0cae802d",
  1560 => x"8e8d2d02",
  1561 => x"84050d04",
  1562 => x"02fc050d",
  1563 => x"725170fd",
  1564 => x"2ead3870",
  1565 => x"fd248a38",
  1566 => x"70fc2e80",
  1567 => x"c438b1c9",
  1568 => x"0470fe2e",
  1569 => x"b13870ff",
  1570 => x"2e098106",
  1571 => x"bc38b98c",
  1572 => x"08517080",
  1573 => x"2eb338ff",
  1574 => x"11b98c0c",
  1575 => x"b1c904b9",
  1576 => x"8c08f005",
  1577 => x"70b98c0c",
  1578 => x"51708025",
  1579 => x"9c38800b",
  1580 => x"b98c0cb1",
  1581 => x"c904b98c",
  1582 => x"088105b9",
  1583 => x"8c0cb1c9",
  1584 => x"04b98c08",
  1585 => x"9005b98c",
  1586 => x"0cae802d",
  1587 => x"8e8d2d02",
  1588 => x"84050d04",
  1589 => x"02fc050d",
  1590 => x"800bb98c",
  1591 => x"0cae802d",
  1592 => x"8d912db9",
  1593 => x"9008b8fc",
  1594 => x"0cb7d851",
  1595 => x"8fa82d02",
  1596 => x"84050d04",
  1597 => x"7180c0c0",
  1598 => x"0c040000",
  1599 => x"00ffffff",
  1600 => x"ff00ffff",
  1601 => x"ffff00ff",
  1602 => x"ffffff00",
  1603 => x"52657365",
  1604 => x"74000000",
  1605 => x"52474220",
  1606 => x"5363616c",
  1607 => x"696e6720",
  1608 => x"10000000",
  1609 => x"5363616e",
  1610 => x"6c696e65",
  1611 => x"73000000",
  1612 => x"416e696d",
  1613 => x"61746500",
  1614 => x"4c6f6164",
  1615 => x"20696d61",
  1616 => x"67652010",
  1617 => x"00000000",
  1618 => x"45786974",
  1619 => x"00000000",
  1620 => x"54657374",
  1621 => x"20706174",
  1622 => x"7465726e",
  1623 => x"20310000",
  1624 => x"54657374",
  1625 => x"20706174",
  1626 => x"7465726e",
  1627 => x"20320000",
  1628 => x"54657374",
  1629 => x"20706174",
  1630 => x"7465726e",
  1631 => x"20330000",
  1632 => x"54657374",
  1633 => x"20706174",
  1634 => x"7465726e",
  1635 => x"20340000",
  1636 => x"52656400",
  1637 => x"47726565",
  1638 => x"6e000000",
  1639 => x"426c7565",
  1640 => x"00000000",
  1641 => x"496e6974",
  1642 => x"69616c20",
  1643 => x"524f4d20",
  1644 => x"6c6f6164",
  1645 => x"696e6720",
  1646 => x"6661696c",
  1647 => x"65640000",
  1648 => x"4f4b0000",
  1649 => x"496e6974",
  1650 => x"69616c69",
  1651 => x"7a696e67",
  1652 => x"20534420",
  1653 => x"63617264",
  1654 => x"0a000000",
  1655 => x"4c6f6164",
  1656 => x"696e6720",
  1657 => x"696e6974",
  1658 => x"69616c20",
  1659 => x"524f4d2e",
  1660 => x"2e2e0a00",
  1661 => x"50494331",
  1662 => x"20202020",
  1663 => x"52415700",
  1664 => x"16200000",
  1665 => x"14200000",
  1666 => x"15200000",
  1667 => x"53442069",
  1668 => x"6e69742e",
  1669 => x"2e2e0a00",
  1670 => x"53442063",
  1671 => x"61726420",
  1672 => x"72657365",
  1673 => x"74206661",
  1674 => x"696c6564",
  1675 => x"210a0000",
  1676 => x"53444843",
  1677 => x"20657272",
  1678 => x"6f72210a",
  1679 => x"00000000",
  1680 => x"57726974",
  1681 => x"65206661",
  1682 => x"696c6564",
  1683 => x"0a000000",
  1684 => x"52656164",
  1685 => x"20666169",
  1686 => x"6c65640a",
  1687 => x"00000000",
  1688 => x"43617264",
  1689 => x"20696e69",
  1690 => x"74206661",
  1691 => x"696c6564",
  1692 => x"0a000000",
  1693 => x"46415431",
  1694 => x"36202020",
  1695 => x"00000000",
  1696 => x"46415433",
  1697 => x"32202020",
  1698 => x"00000000",
  1699 => x"4e6f2070",
  1700 => x"61727469",
  1701 => x"74696f6e",
  1702 => x"20736967",
  1703 => x"0a000000",
  1704 => x"42616420",
  1705 => x"70617274",
  1706 => x"0a000000",
  1707 => x"4261636b",
  1708 => x"00000000",
  1709 => x"00000002",
  1710 => x"00000002",
  1711 => x"0000190c",
  1712 => x"00000352",
  1713 => x"00000003",
  1714 => x"00001b18",
  1715 => x"00000004",
  1716 => x"00000004",
  1717 => x"00001914",
  1718 => x"00001b28",
  1719 => x"00000001",
  1720 => x"00001924",
  1721 => x"00000000",
  1722 => x"00000002",
  1723 => x"00001930",
  1724 => x"00000324",
  1725 => x"00000002",
  1726 => x"00001938",
  1727 => x"000018d4",
  1728 => x"00000002",
  1729 => x"00001948",
  1730 => x"000006ab",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00001950",
  1735 => x"00001960",
  1736 => x"00001970",
  1737 => x"00001980",
  1738 => x"00000005",
  1739 => x"00001990",
  1740 => x"00000010",
  1741 => x"00000005",
  1742 => x"00001994",
  1743 => x"00000010",
  1744 => x"00000005",
  1745 => x"0000199c",
  1746 => x"00000010",
  1747 => x"00000004",
  1748 => x"00001948",
  1749 => x"00001ab8",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000004",
  1754 => x"000019a4",
  1755 => x"00001b64",
  1756 => x"00000004",
  1757 => x"000019c0",
  1758 => x"00001ab8",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000002",
  1783 => x"00002044",
  1784 => x"000016cd",
  1785 => x"00000002",
  1786 => x"00002062",
  1787 => x"000016cd",
  1788 => x"00000002",
  1789 => x"00002080",
  1790 => x"000016cd",
  1791 => x"00000002",
  1792 => x"0000209e",
  1793 => x"000016cd",
  1794 => x"00000002",
  1795 => x"000020bc",
  1796 => x"000016cd",
  1797 => x"00000002",
  1798 => x"000020da",
  1799 => x"000016cd",
  1800 => x"00000002",
  1801 => x"000020f8",
  1802 => x"000016cd",
  1803 => x"00000002",
  1804 => x"00002116",
  1805 => x"000016cd",
  1806 => x"00000002",
  1807 => x"00002134",
  1808 => x"000016cd",
  1809 => x"00000002",
  1810 => x"00002152",
  1811 => x"000016cd",
  1812 => x"00000002",
  1813 => x"00002170",
  1814 => x"000016cd",
  1815 => x"00000002",
  1816 => x"0000218e",
  1817 => x"000016cd",
  1818 => x"00000002",
  1819 => x"000021ac",
  1820 => x"000016cd",
  1821 => x"00000004",
  1822 => x"00001aac",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00001868",
  1827 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

